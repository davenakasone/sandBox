/*
    the hello-world of verilog
*/

module hello(A,B);
    input A;
    output B;
    assign B = A;
endmodule

////////~~~~~~~~END>  hello.v

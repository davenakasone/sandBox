/*
    showing JAL on FPGA
*/

`timescale 1ns/1ns
`define HALF 5         // half cycle, time between posedge and negedge
`define NANO_SPIN 0    // reps until last instruction
`define SAFETY 15      // kill after this many of instructions, stops oo loop                                       

// original "testbench.v"  ,  file 1 of 16
////~~~~
/*
    should be updated to reflect instruction sets
    control the MACROS for selecting the proper instructions to test
    only makes DUT from top module, 
        member access to see internals, or turn on individual DEBUG macros
*/
module test_bench();
    reg clock;
    reg reset;
    wire [6:0] lsb_reg;
    wire memwrite;
    wire ready;

    powerTop DUT (
                    .clk(clock),
                    .reset(reset),
                    .lsb_reg(lsb_reg),
                    .memwrite(memwrite),
                    .ready(ready)
                );

    reg printing;
    integer idx;
    reg sim_success;
    integer play_time;
    reg access_complete;

    initial begin
        printing = 1'b0;
        idx = 1;
        sim_success = 1'b0;
        access_complete = 1'b0;
        play_time = `NANO_SPIN;  // change in macro

        reset <= 1; 
        # `HALF; 
        # `HALF; 
        reset <= 0;
        # 2;
        printing = 1'b1;

        $write("\n testing verison:  \"jal\"  with sub-routine ,");
        $write("  success means M[0x50] = 0xA\n");
    end

    always begin
        clock <= 1'b0;
        # `HALF; 
        clock <= 1'b1;
        # `HALF; 
    end

    // instructions in  "jal_test.dat"  ,  success means M[80] = 10
    always @ (negedge clock) begin
        if (memwrite == 1'b1 && ready == 1'b1 && lsb_reg == 7'b0001000) begin 
            sim_success = 1'b1;
            access_complete = 1'b1;
        end
        else begin
            sim_success = 1'b0;
        end
    end

    always @ (negedge clock) begin
        #1;
        if (printing) begin
            idx = idx + 1;
        end

        play_time = (access_complete == 1'b1) ? play_time - 1 : play_time;

        if (play_time < 0 || idx > `SAFETY) begin
            if (sim_success == 1'b1) begin
                $write("\n\n\tSimulation SUCCESS\n");
            end
            else begin
                $write("\n\n\tSimulation FAIL\n");
            end
            $write("\n\n\t\t ~ ~ ~ TEST COMPLETE ~ ~ ~    %9t ns\n\n", $time);
            $finish;
        end 
    end

endmodule


////~~~~ for the FPGA
module powerTop (
                    input wire clk,
                    input wire reset,
                    output reg [6:0] lsb_reg,
                    output wire memwrite,
                    output reg ready
                );

    wire [31:0] writedata;
    wire [31:0] dataadr;
    wire [6:0] catch;

    m_main inst_top (
                    .clock(clk),
                    .reset(reset),
                    .writedata(writedata),
                    .dataadr(dataadr),
                    .memwrite(memwrite)
                );
    
    seg7_dig1 get_dig (
                        .cntl(writedata[3:0]),
                        .disp(catch)
                    );
    
    always @ (*) begin
        if (memwrite == 1'b1) begin
            if (dataadr === 80 & writedata === 10) begin
                ready <= 1'b1;
                lsb_reg <= catch;
            end 
        end
        else begin
            ready <= 1'b0;
            lsb_reg <= 7'b1111_111;
        end
        
    end
    
endmodule


////~~~~
module seg7_dig1(
                input [3:0] cntl,
                output reg [6:0] disp
            );

    parameter ON = 1'b0;
    parameter OFF = 1'b1;

    always @ (*) begin
        disp = {7{OFF}};
        case (cntl)
            4'b0000 : disp[5:0] = {6{ON}};
            4'b0001 : disp[2:1] = {2{ON}};
            4'b0010 :
                begin
                    disp[1:0] = {2{ON}};
                    disp[6] = ON;
                    disp[4:3] = {2{ON}};
                end
            4'b0011 :
                begin
                    disp[3:0] = {4{ON}};
                    disp[6] = ON;
                end
            4'b0100 :
                begin
                    disp[2:1] = {2{ON}};
                    disp[6:5] = {2{ON}};
                end 
            4'b0101 :
                begin
                    disp[0] = ON;
                    disp[3:2] = {2{ON}};
                    disp[6:5] = {2{ON}};
                end
            4'b0110 :
                begin
                    disp[0] = ON;
                    disp[6:2] = {5{ON}};
                end
            4'b0111 : disp[2:0] = {3{ON}};
            4'b1000 : disp[6:0] = {7{ON}};
            4'b1001 :
                begin
                    disp[6:0] = {7{ON}};
                    disp[4:3] = {2{OFF}};
                end
            4'b1010 :
                begin
                    disp = {7{ON}};
                    disp[3] = OFF;
                end
            default : disp = {7{OFF}};
        endcase
    end
endmodule


// original "top.v"  ,  file 2 of 16
////~~~~
/*
    the applied microprocessor
    combines: instruction_memory, dynamic_memory, and mips
    module that should be tested, not a diagram component
*/
module m_main (
                input wire clock, 
                input wire reset,
                output wire [31:0] writedata, 
                output wire [31:0] dataadr,
                output wire memwrite
            );

    wire [31:0] pc;
    wire [31:0] instr; 
    wire [31:0] readdata;

    mips_dp_cu mips (clock, reset, pc, instr, memwrite, dataadr, writedata, readdata);
    instruction_memory imem (pc[7:2], instr);
    dynamic_memory dmem (clock, memwrite, dataadr, writedata, readdata);

endmodule


// original "mips.v"  ,  file 3 of 16
////~~~~
/*
    mips has 4 fundamental units: 
        program counter, instruction memory, register file, and data memory
    this module only combines the control unit and data path
    be careful for those originally missing wires (see comments)
        verify with:
            DEBUG_mips_dp_cu
*/
module mips_dp_cu (
                    input wire clock, 
                    input wire reset,
                    output wire [31:0] pc,
                    input wire [31:0] instr,
                    output wire memwrite,
                    output wire [31:0] aluout, 
                    output wire [31:0] writedata,
                    input wire [31:0] readdata
                );

    wire memtoreg;
    wire alusrc;
    wire regdst;
    wire regwrite;
    wire jump;
    wire [2:0] alucontrol;
    wire zero;     
    wire pcsrc;    
    wire sig_ori;  
    wire sig_jr;   
    wire sig_lui;
    wire sig_jal;

    control_unit CU (
                    .op(instr[31:26]), 
                    .funct(instr[5:0]),
                    .zero(zero),
                    .memtoreg(memtoreg), 
                    .memwrite(memwrite),
                    .pcsrc(pcsrc), 
                    .alusrc(alusrc),
                    .regdst(regdst), 
                    .regwrite(regwrite),
                    .jump(jump),
                    .sig_ori(sig_ori),  
                    .sig_jr(sig_jr),    
                    .sig_lui(sig_lui), 
                    .sig_jal(sig_jal), 
                    .alucontrol(alucontrol)
                );
    
    data_path DP (
                    .clock(clock), 
                    .reset(reset),
                    .memtoreg(memtoreg), 
                    .pcsrc(pcsrc),
                    .alusrc(alusrc), 
                    .regdst(regdst),
                    .regwrite(regwrite), 
                    .jump(jump),
                    .sig_ori(sig_ori),  
                    .sig_jr(sig_jr),    
                    .sig_lui(sig_lui), 
                    .sig_jal(sig_jal), 
                    .alucontrol(alucontrol),
                    .zero(zero),
                    .pc(pc),
                    .instr(instr),
                    .aluout(aluout), 
                    .writedata(writedata),
                    .readdata(readdata)
                );
endmodule


// original "imem.v"  ,  file 4 of 16
////~~~~
/*
    instruction memory wouldn't really be a ROM
    drive instructions from intially reading a file
    verify with:
        DEBUG_INITIAL
        BASE_TEST_1
        BASE_TEST_2
        ORI_TEST
        JR_TEST
        SLLV_LUI_TEST
        DEBUG_instruction_memory
*/
module instruction_memory (
                                input wire [5:0] a, 
                                output wire [31:0] rd
                            );

    reg [31:0] RAM[63:0];  // limited memory

    `ifdef DEBUG_INITIAL
        reg [31:0] temp;
        integer ii;
    `endif
    
    initial begin
        RAM[0] = 32'h2004_0002;
        RAM[1] = 32'h2005_0003;
        RAM[2] = 32'h0C00_0005;
        RAM[3] = 32'h0800_0009;
        RAM[4] = 32'h2010_0001;
        RAM[5] = 32'h0085_4020;
        RAM[6] = 32'h2009_0001;
        RAM[7] = 32'h0128_1004;
        RAM[8] = 32'h03E0_0008;
        RAM[9] = 32'hAC02_0050;
    end

    assign rd = RAM[a];  // word aligned, always reads to output

endmodule


// original "dmem.v"  ,  file 5 of 16
////~~~~
/*
    data memory reads in combination
    writes synchronously on positive edge of clock
    verify with:
        DEBUG_dynamic_memory
*/
module dynamic_memory (
                input wire clock, 
                input wire we,
                input wire [31:0] a, 
                input wire [31:0] wd,
                output [31:0] rd
            );

    reg [31:0] RAM[63:0];

    assign rd = RAM[a[31:2]]; // word aligned

    always @ (posedge clock) begin
        if (we) RAM[a[31:2]] <= wd;
    end

endmodule


// original "controller.v"  ,  file 6 of 16
////~~~~
/*
    sub-components of ALU decoder and main decoder
    implies AND gate for pcsrc
    update as instruction set changes
*/
module control_unit (
                    input wire [5:0] op, 
                    input wire [5:0] funct,
                    input wire zero,
                    output wire memtoreg, 
                    output wire memwrite,
                    output wire pcsrc, 
                    output wire alusrc,
                    output wire regdst, 
                    output wire regwrite,
                    output wire jump,
                    output wire sig_ori,  
                    output wire sig_jr,   
                    output wire sig_lui, 
                    output wire sig_jal, 
                    output wire [2:0] alucontrol
                );

    wire [1:0] aluop;
    wire branch;

    maindec MD (
                    .op(op), 
                    .funct(funct),
                    .memtoreg(memtoreg), 
                    .memwrite(memwrite), 
                    .branch(branch), 
                    .alusrc(alusrc),
                    .regdst(regdst), 
                    .regwrite(regwrite), 
                    .jump(jump), 
                    .sig_ori(sig_ori),  
                    .sig_jr(sig_jr),    
                    .sig_lui(sig_lui),
                    .sig_jal(sig_jal),  
                    .aluop(aluop)
                );

    aludec AD (funct, aluop, alucontrol);

    assign pcsrc = branch & zero;  // the AND gate in diagram

endmodule


// original "maindec.v"  ,  file 7 of 16
////~~~~
/*
    takes opcode and produces control signals except branch
    branching is done by controller module as an outside logic
    checks the opcode and produces 9 control signals {control word table}
*/
module maindec (
                    input wire [5:0] op, 
                    input wire [5:0] funct,
                    output wire memtoreg, 
                    output wire memwrite, 
                    output wire branch, 
                    output wire alusrc,
                    output wire regdst, 
                    output wire regwrite, 
                    output wire jump, 
                    output wire sig_ori,  
                    output wire sig_jr,   
                    output wire sig_lui,  
                    output wire sig_jal,
                    output wire [1:0] aluop
                );

    reg [12:0] controls; 

    assign {regwrite, regdst, alusrc, branch, memwrite, memtoreg, 
        aluop, jump, sig_ori, sig_jr, sig_lui, sig_jal} = controls; 

    always @ (*) begin // new
        case(op)
            6'b000_000 :                                       
                        begin
                            if (funct == 6'b001_000) begin
                                controls <= 13'b0_0_0_0_0_0_10_0_0_1_0_0; // R-type, is JR
                            end
                            else begin
                               controls <= 13'b1_1_0_0_0_0_10_0_0_0_0_0; // R-type, not jr 
                            end   
                        end
            6'b100_011 :  controls <= 13'b1_0_1_0_0_1_00_0_0_0_0_0;    // lw
            6'b101_011 :  controls <= 13'b0_0_1_0_1_0_00_0_0_0_0_0;    // sw
            6'b000_100 :  controls <= 13'b0_0_0_1_0_0_01_0_0_0_0_0;    // beq
            6'b001_000 :  controls <= 13'b1_0_1_0_0_0_00_0_0_0_0_0;    // addi
            6'b000_010 :  controls <= 13'b0_0_0_0_0_0_00_1_0_0_0_0;    // j
            6'b001_101 :  controls <= 13'b1_0_1_0_0_0_11_0_1_0_0_0;    // ori
            6'b001_111 :  controls <= 13'b1_0_0_0_0_0_00_0_0_0_1_0;    // lui
            6'b000_011 :  controls <= 13'b1_0_0_0_0_0_00_1_0_0_0_1;    // jal
            default    :  controls <= 13'bX_X_X_X_X_X_XX_X_X_X_X_X;    // any
        endcase
    end

endmodule


// original "aludec.v"  ,  file 8 of 16
////~~~~
/*
    this will get overloaded quickly if more signals are needed
*/
module aludec (
                    input wire [5:0] funct,
                    input wire [1:0] aluop,
                    output reg [2:0] alucontrol
            );

    always @ (*) begin
        if (aluop == 2'b00) begin
            alucontrol <= 3'b010; // add
        end
        else if (aluop == 2'b01) begin
            alucontrol <= 3'b110; // sub
        end
        else if (aluop == 2'b11) begin
            alucontrol <= 3'b001; // if more than "ori" use 2'b11, make case statement
        end
        else begin // R-type  2'b10 case
            case(funct) 
                6'b100_000 : alucontrol <= 3'b010; // add
                6'b100_010 : alucontrol <= 3'b110; // sub
                6'b100_100 : alucontrol <= 3'b000; // and
                6'b100_101 : alucontrol <= 3'b001; // or
                6'b101_010 : alucontrol <= 3'b111; // slt
                6'b000_100 : alucontrol <= 3'b101; // sllv
                default    : alucontrol <= 3'bxxx; // catch all {jr}
            endcase
        end
    end

endmodule


// original "datapth.v"  ,  file 9 of 16
////~~~~
/*
    control signals determine operation
    the data path and control unit work together as usual
*/
module data_path (
                    input wire clock, 
                    input wire reset,
                    input wire memtoreg, 
                    input wire pcsrc,
                    input wire alusrc, 
                    input wire regdst,
                    input wire regwrite, 
                    input wire jump,
                    input wire sig_ori,  
                    input wire sig_jr,   
                    input wire sig_lui, 
                    input wire sig_jal,
                    input wire [2:0] alucontrol,
                    output wire zero,
                    output wire [31:0] pc,
                    input wire [31:0] instr,
                    output wire [31:0] aluout, 
                    output wire [31:0] writedata,
                    input wire [31:0] readdata
                );

    wire [4:0] writereg;
    wire [31:0] pcnext;
    wire [31:0] pcnextbr;
    wire [31:0] pcplus4;
    wire [31:0] pcbranch;
    wire [31:0] signimm;
    wire [31:0] signimmsh;
    wire [31:0] srca;
    wire [31:0] srcb;
    wire [31:0] result;
    wire [31:0] zeroXimm;        
    wire [31:0] extend_mux_out;  
    wire [31:0] jr_mux_out;      
    wire [31:0] write_to_rf;      
    wire [31:0] zero_full;   
    wire [4:0] from_wrmux;  
    wire [31:0] from_lui_mux;   

    // next PC logic
    program_counter #(32) pcreg (clock, reset, pcnext, pc);
    adder pcadd1 (pc, 32'b100, pcplus4);
    shift_left_2 immsh (signimm, signimmsh); 
    adder pcadd2 (pcplus4, signimmsh, pcbranch);
    mux_2_to_1 #(32) pcbrmux (pcplus4, pcbranch, pcsrc, pcnextbr);
    mux_2_to_1 #(32) jr_mux (pcnextbr, srca, sig_jr, jr_mux_out); 
    mux_2_to_1 #(32) pcmux (jr_mux_out, {pcplus4[31:28], instr[25:0], 2'b00}, jump, pcnext); 

    // register file logic
    register_file RF (clock, regwrite, instr[25:21], instr[20:16], writereg, write_to_rf, srca, writedata); 
    mux_2_to_1 #(5) wrmux (instr[20:16], instr[15:11], regdst, from_wrmux);
    mux_2_to_1 #(5) wrmux_jal (from_wrmux, 5'b11111, sig_jal, writereg);
    mux_2_to_1 #(32) resmux (aluout, readdata, memtoreg, result);
    mux_2_to_1 #(32) lui_mux (result, zero_full, sig_lui, from_lui_mux); 
    mux_2_to_1 #(32) mux_rf_write(from_lui_mux, pcplus4, sig_jal, write_to_rf);
    sign_extend SE (instr[15:0], signimm);
    zero_extend ZE (instr[15:0], zeroXimm);  
    zero_filler ZF (instr[15:0], zero_full);  

    // ALU logic
    mux_2_to_1 #(32) srcbmux (writedata, extend_mux_out, alusrc, srcb); 
    mux_2_to_1 #(32) extend_mux (signimm, zeroXimm, sig_ori, extend_mux_out);  
    alu ALU (srca, srcb, alucontrol, aluout, zero);

endmodule


// original "flopr.v"  ,  file 10 of 16
////~~~~
/*
    32 D flip-flops to represent the program counter
    notice it resets to 8'h0000_0000  (change as needed)
*/
module program_counter # (parameter WIDTH = 8) (
                                        input wire clock, 
                                        input wire reset,
                                        input wire [WIDTH-1:0] d,
                                        output reg [WIDTH-1:0] q
                                    );

    always @ (posedge clock or posedge reset) begin
        q <= (reset) ? 0 : d;
    end

endmodule


// original "adder.v"  ,  file 11 of 16
////~~~~
/*
    there is not much going on here
    be careful for overflow
*/
module adder (
                input wire [31:0] a, 
                input wire [31:0] b, 
                output wire [31:0] y
            );

    assign y = a + b;

endmodule


// original "sl2.v"  ,  file 12 of 16
////~~~~
/*
    appends two zeros from the right of LSB 
    for 26-bit immediate field provided as input
    shift left by 2 bits uses concatenation
        26 + 2 = 28 bits out [27:0]
*/
module shift_left_2 (
                input wire [31:0] a, 
                output wire [31:0] y
            );

    assign y = {a[25:0], 2'b00};

endmodule


// original "mux2.v"  ,  file 13 of 16
////~~~~
/*
    ordinary 2:1 MUX using parameterized inputs
    Please note, it is limited to 8 as both 
    addresses for instruction and data memory are limited to 6.
    data in the test code are in the range 0-255
    For the real design the width is 8
*/ 
module mux_2_to_1 # (parameter WIDTH = 8) (
                                        input wire [WIDTH-1:0] d0, 
                                        input wire [WIDTH-1:0] d1, 
                                        input wire s,
                                        output wire [WIDTH-1:0] y
                                    );

    assign y = (s) ? d1 : d0;

endmodule


// original "regfile.v"  ,  file 14 of 16
////~~~~
/*
    this is one of the fundamental elements of the CPU
    3-ported register file
    it reads 2 ports out in combination, 
    but writes sychrousnously (posedge)
    register 0 hardwired to 0
*/
module register_file (
                        input wire clock, 
                        input wire we3,
                        input wire [4:0] ra1, 
                        input wire [4:0] ra2, 
                        input wire [4:0] wa3,
                        input wire [31:0] wd3,
                        output wire [31:0] rd1, 
                        output wire [31:0]rd2
                    );

    reg [31:0] rf[31:0];
    
    always @ (posedge clock) begin
        if (we3) rf[wa3] <= wd3;
    end

    // notice the effective hard-wire rf[0] = 0
    assign rd1 = (ra1 != 0) ? rf[ra1] : 0; 
    assign rd2 = (ra2 != 0) ? rf[ra2] : 0; 

endmodule


// original "signext.v"  ,  file 15 of 16
////~~~~
/*
    effective sign externsion 
    concatenates to output a 32-bit number
    copies the 16th bit of input "a[15]"  
        to upper of output "y[31:16]"
*/
module sign_extend (
                    input wire [15:0] a,
                    output wire [31:0] y
                );

    assign y = {{16{a[15]}}, a};

endmodule


// original "alu.v"  ,  file 16 of 16
////~~~~
/*
    ordinary ALU that also outputs zero flag
    it still has room to add more
*/
module alu (
                input wire [31:0] a,
                input wire [31:0] b,
                input wire [2:0] sel, 
                output reg [31:0] out, 
                output reg zero
            );
  
    initial begin
        out = 0;
        zero =1'b0;
    end
    
    always @ (*) begin 
        case(sel) 
            3'b000 : 
	            begin
		            out = a & b; 
		            if (out == 0) zero = 1;  
		            else zero = 0;
                end                   
            3'b001 :
	            begin
		            out= a | b; 
		            if (out == 0) zero = 1;  
		            else zero = 0; 
                end	
            3'b010 : 
	            begin
		            out = a + b;  
		            if (out == 0) zero = 1;  
                    else zero = 0;
                end  
            3'b101 : 
	            begin
		            out = b << a;
                end  	
            3'b110 : 
	            begin
		            out = a - b;  
		            if (out == 0) zero = 1;  
		            else zero = 0;
                end              
            3'b111 : 
                begin
		            if ( a < b) out = 1;  
		            else out = 0;
                end 
            default : 
                begin
                    out = 0;
                    zero = 0;
                end
        endcase
    end

endmodule


////~~~~
/*
    zero extends the immidate 
    from 16-bits to 32-bits by concatenation
*/
module zero_extend (
                    input wire [15:0] a,
                    output wire [31:0] y
                );

    assign y = {16'h0000, a};

endmodule


////~~~~
/*
    zero fills LSBs after immidate 
    {immediate, 16{0}}
*/
module zero_filler (
                    input wire [15:0] a,
                    output wire [31:0] y
                );

    assign y = {a,16'h0000};

endmodule


////////~~~~~~~~END>  mips_single_enhanced.v
